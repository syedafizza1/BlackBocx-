module orGate(output Y, input A, B);
   or(Y, A, B); 
endmodule